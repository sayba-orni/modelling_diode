* C:\Users\Lenovo\3D Objects\DIODE_FINAL_PROJECT\Diode\Schematic2.sch

* Schematics Version 9.2
* Wed Mar 01 13:43:45 2023



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "Schematic2.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
