* C:\Users\Lenovo\3D Objects\DIODE_FINAL_PROJECT\Diode\2.sch

* Schematics Version 9.2
* Wed Mar 01 08:43:44 2023



** Analysis setup **
.OP 
.LIB "C:\Users\USER\Desktop\Schematic1.lib"


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "2.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
